module Lab7part1

endmodule
